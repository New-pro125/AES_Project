module shiftRows_tb;
reg [127:0] din;
wire [127:0] dout;
initial 
begin
        din=128'hd42711aee0bf98f1b8b45de51e415230;
end
shiftRows u (.din(din),.dout(dout));
endmodule