
module INVshiftRows_tb;
reg [127:0] din;
wire [127:0] dout;
initial 
begin
        din=128'hd4bf5d30e0b452aeb84111f11e2798e5;
end
invShiftRows u (.din(din),.dout(dout));
endmodule